--
-- Copyright (c) 2018, UPC
-- All rights reserved.
-- 

library ieee;
use ieee.std_logic_1164.all;

package retardos_bcd_pkg is

constant retsumbin: time := 2 ns;
constant retmayor9: time := 1 ns;
constant rets1bit: time := 1 ns;
constant retc9: time := 1 ns;
constant retmux: time := 1 ns;
constant retBCDaDPD: time := 1 ns;
constant retDPDaBCD: time := 1 ns;

end package retardos_bcd_pkg;

